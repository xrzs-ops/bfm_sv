module uart(
    input   rx,
    output  tx
);

    assign tx = rx;
    
endmodule